`define MASTER_NUM      2
`define SLAVE_NUM       8
`define W_ID_LEN        4
`define R_ID_LEN        4
`define EXTRA_ID_LEN    1
`define ADDR_WIDTH      32
`define DATA_WIDTH      64
`define W_BUF_DEPTH     3
`define R_BUF_DEPTH     3